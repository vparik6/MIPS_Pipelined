/*
mipscpu_tb.sv
*/

module mipscpu_tb.sv


endmodule