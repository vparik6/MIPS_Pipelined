/*
mux.sv
-consider reusability (with parameter)
*/


module mux_pc

endmodule


module mux_ex1


endmodule



module mux_ex1


endmodule



module mux_wb


endmodule