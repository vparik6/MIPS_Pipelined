/*
StallUnit.sv
input:
output:
*/

module StallUnit

endmodule