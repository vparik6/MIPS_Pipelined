/*
ProgramCounter.sv
input:clk,reset,pc_in,stallF
output:pc_out
*/

module ProgramCounter



endmodule