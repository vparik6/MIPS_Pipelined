/*
DataMemory.sv
input: clk,MemWriteM,ALUOutM,WriteDataM
output: ReadDataM
*/

module DataMemory

endmodule