/*
MEM_WB.sv
input: clk,reset,RegWriteM,MemtoRegM,ReadDataM,ALUOutM,WriteRegM
output: RegWriteW,MemtoRegW,ReadDataW,ALUOutW,WriteRegW
*/ 

module MEM_WB

endmodule