/*
ID_EX.sv
input: clk,reset,FlushE,RegWriteD,MemtoRegD,MemWriteD,ALUControlD,ALUSrcD,RegDstD,BranchD,rd1_ID,rd2_ID,RsD,RtD,RdD,SignImmD,PCPlus4D
output: rd1_EX,rd2_EX,RsE,RtE,RdE,SignImmE,PCPlus4E
*/

module ID_EX

endmodule