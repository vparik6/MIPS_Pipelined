/*
IF_ID.sv
input: clk,reset,InstrF,PCPlus4F,stallD
output: InstrD,PCPlus4D
*/

module IF_ID.sv

endmodule