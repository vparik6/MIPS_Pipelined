/*
ControlUnit.sv
input: InstrD[31:26],InstrD[5:0]
output: RegWriteD,MemtoRegD,MemWriteD,ALUControlD,ALUSrcD,RegDstD,BranchD
*/

module ControlUnit

endmodule