/*
alu.sv
input: ALUControlE,SrcAE,SrcBE
output: ZeroE,ALUOutE
*/

module alu

endmodule