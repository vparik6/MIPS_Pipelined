/*
InstructionMemory.sv
input: pc_out
output: InstrF
*/

module InstructionMemory

endmodule